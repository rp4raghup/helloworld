module helloworld;
initial $display("hello world");
endmodule
